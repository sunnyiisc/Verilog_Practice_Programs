module hello_world;
    initial begin
        $display("Hello Supantha");
        #10 $finish;
    end
endmodule